-- Create Date:    18:21:15 07/12/2022 
-- Design Name: 
-- Module Name:    SistemaSecuencial - Behavioral 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SistemaSecuencial is
end SistemaSecuencial;

architecture Behavioral of SistemaSecuencial is

begin


end Behavioral;

