-- Create Date:    18:19:23 07/12/2022 
-- Design Name: 
-- Module Name:    DetectorSecuencia - Behavioral 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DetectorSecuencia is
end DetectorSecuencia;

architecture Behavioral of DetectorSecuencia is

begin


end Behavioral;

